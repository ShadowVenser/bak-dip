[info] welcome to sbt 1.10.7 (Temurin Java 1.8.0_442)
[info] loading project definition from /home/venser/bak-dip/chisel/testings/example/project
[info] loading settings for project root from build.sbt...
[info] set current project to %NAME% (in build file:/home/venser/bak-dip/chisel/testings/example/)
[info] compiling 1 Scala source to /home/venser/bak-dip/chisel/testings/example/target/scala-2.13/classes ...
[info] done compiling
[info] compiling 1 Scala source to /home/venser/bak-dip/chisel/testings/example/target/scala-2.13/classes ...
[info] done compiling
[info] running Main 
// Generated by CIRCT firtool-1.114.1
module NandGate(
  input  x1,
         x2,
  output y
);

  assign y = ~(x1 & x2);
endmodule


// ----- 8< ----- FILE "verification/cover/layers-NandGate-Verification-Cover.sv" ----- 8< -----

// Generated by CIRCT firtool-1.114.1
`include "verification/layers-NandGate-Verification.sv"
`ifndef layers_NandGate_Verification_Cover
`define layers_NandGate_Verification_Cover
`endif // layers_NandGate_Verification_Cover

// ----- 8< ----- FILE "verification/assume/layers-NandGate-Verification-Assume.sv" ----- 8< -----

// Generated by CIRCT firtool-1.114.1
`include "verification/layers-NandGate-Verification.sv"
`ifndef layers_NandGate_Verification_Assume
`define layers_NandGate_Verification_Assume
`endif // layers_NandGate_Verification_Assume

// ----- 8< ----- FILE "verification/assert/layers-NandGate-Verification-Assert.sv" ----- 8< -----

// Generated by CIRCT firtool-1.114.1
`include "verification/layers-NandGate-Verification.sv"
`ifndef layers_NandGate_Verification_Assert
`define layers_NandGate_Verification_Assert
`endif // layers_NandGate_Verification_Assert

// ----- 8< ----- FILE "verification/layers-NandGate-Verification.sv" ----- 8< -----

// Generated by CIRCT firtool-1.114.1
`ifndef layers_NandGate_Verification
`define layers_NandGate_Verification
`endif // layers_NandGate_Verification

// Generated by CIRCT firtool-1.114.1
module SyncMux(
  input         clk,
                clr_n,
  input  [15:0] x1,
                x2,
  input         addr,
  output [15:0] y
);

  wire        _asyncReset_T = ~clr_n;
  reg  [15:0] y_reg;
  always @(posedge clk or posedge _asyncReset_T) begin
    if (_asyncReset_T)
      y_reg <= 16'h0;
    else
      y_reg <= addr ? x2 : x1;
  end // always @(posedge, posedge)
  `ifdef ENABLE_INITIAL_REG_
    `ifdef FIRRTL_BEFORE_INITIAL
      `FIRRTL_BEFORE_INITIAL
    `endif // FIRRTL_BEFORE_INITIAL
    initial begin
      if (_asyncReset_T)
        y_reg = 16'h0;
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL
      `FIRRTL_AFTER_INITIAL
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  assign y = y_reg;
endmodule


// ----- 8< ----- FILE "verification/cover/layers-SyncMux-Verification-Cover.sv" ----- 8< -----

// Generated by CIRCT firtool-1.114.1
`include "verification/layers-SyncMux-Verification.sv"
`ifndef layers_SyncMux_Verification_Cover
`define layers_SyncMux_Verification_Cover
`endif // layers_SyncMux_Verification_Cover

// ----- 8< ----- FILE "verification/assume/layers-SyncMux-Verification-Assume.sv" ----- 8< -----

// Generated by CIRCT firtool-1.114.1
`include "verification/layers-SyncMux-Verification.sv"
`ifndef layers_SyncMux_Verification_Assume
`define layers_SyncMux_Verification_Assume
`endif // layers_SyncMux_Verification_Assume

// ----- 8< ----- FILE "verification/assert/layers-SyncMux-Verification-Assert.sv" ----- 8< -----

// Generated by CIRCT firtool-1.114.1
`include "verification/layers-SyncMux-Verification.sv"
`ifndef layers_SyncMux_Verification_Assert
`define layers_SyncMux_Verification_Assert
`endif // layers_SyncMux_Verification_Assert

// ----- 8< ----- FILE "verification/layers-SyncMux-Verification.sv" ----- 8< -----

// Generated by CIRCT firtool-1.114.1
`ifndef layers_SyncMux_Verification
`define layers_SyncMux_Verification
`endif // layers_SyncMux_Verification

[success] Total time: 6 s, completed 22.05.2025 2:48:30
